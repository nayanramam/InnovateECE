module counter_16bit (
    input wire clk,
    input wire rst_n,
    input wire enable,
    output reg [15:0] count
);

always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        count <= 16'h0000;
    end else if (enable) begin
        count <= count + 1'b1;
    end else begin
        count <= count;
    end
end

endmodule